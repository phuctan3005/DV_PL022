package test_pkg;    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import ssp_pkg::*;
    //import env_pkg::*;
    import seq_pkg::*;
    `include "ssp_base_test.sv"
    `include "default_value_test.sv"
endpackage