package ssp_pkg; 
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "ssp_transaction.sv"
    `include "ssp_sequencer.sv"
    `include "ssp_driver.sv"
    `include "ssp_monitor.sv"
    `include "ssp_agent.sv"
    `include "ssp_scoreboard.sv"
    `include "ssp_environment.sv"
endpackage : ssp_pkg