/////////////////////////////