package env_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import ssp_pkg::*;
    `include "ssp_scoreboard.sv"
    `include "ssp_environment.sv"
endpackage